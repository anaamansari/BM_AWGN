`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 03/19/2016 04:08:08 PM
// Design Name: 
// Module Name: LZDfortyeigth
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module LZDfortyeight(
    input [47:0] a,
    output reg [5:0] p,
    output reg v
    );
    
    wire [4:0] p2;
    wire [3:0] p1;
                                                                                                                                                                                                               
   wire v2,v1;
            
            
            LZDthtwo l2(
            .a(a[47:16]),
            .p(p2),
            .v(v2)
            );
            
            LZDsixteen l1(
              .a(a[15:0]),
              .p(p1),
              .v(v1)
            );
            
             always@(a,p1,v1,p2,v2) begin
                            v= v1 | v2;
                             if (v2==0)begin
                              p= {{~v2}, {1'b0,{p1}}};
                              end
                              else begin
                             p= {{~v2}, {p2}};
                              end
                   v <= v1 | v2;
                   end
endmodule
